module Controls_1(
  input [6:0] x,
  input [5:0] y,
  output reg [15:0] oled_data
);

//Define constant as local parameter
//Colour display
localparam GREEN = 16'h07E0;
localparam ORANGE = 16'hFFE0; //Yellow
localparam RED = 16'hF800;
localparam BLACK = 16'h0000;
localparam PURPLE = 16'hF81F;
localparam YELLOW = 16'hFC00;    
localparam BLUE = 16'h001F;
localparam WHITE = 16'hFFFF;
localparam CYAN = 16'hF81F;
localparam MAGENTA = 16'hF81F;
localparam BROWN = 16'h8204;
localparam SKYBLUE = 16'h5FFF;

    //Display Game Control
    wire S1 = ((x >= 20 && x <= 21) && (y >= 5 && y <= 7)) || ((x >= 22 && x <= 23) && (y == 5)) || ((x >= 22 && x <= 23) && (y >= 7 && y <= 9)) || ((x >= 20 && x <= 21) && (y == 9)) ||
              ((x >= 25 && x <= 26) && (y >= 5 && y <= 9)) || ((x >= 27 && x <= 28) && (y == 5)) || ((x == 27) && (y == 7)) || ((x >= 27 && x <= 28) && (y == 9)) ||
              ((x >= 30 && x <= 33) && (y == 5)) || ((x >= 31 && x <= 32) && (y >= 5 && y <= 9)) ||
              ((x >= 35 && x <= 38) && (y == 5)) || ((x >= 36 && x <= 37) && (y >= 5 && y <= 9)) ||
              ((x >= 40 && x <= 43) && (y == 5)) || ((x >= 41 && x <= 42) && (y >= 5 && y <= 9)) || ((x >= 40 && x <= 43) && (y == 9)) ||
              ((x >= 45 && x <= 46) && (y >= 5 && y <= 9)) || ((x == 47) && (y == 5)) || ((x == 48) && (y >= 5 && y <= 9)) ||
              ((x >= 50 && x <= 51) && (y >= 5 && y <= 9)) || ((x >= 52 && x <= 53) && (y == 5)) || ((x == 52) && (y == 9)) || ((x == 53) && (y >= 7 && y <= 9)) ||
                         
              ((x >= 57 && x <= 58) && (y >= 5 && y <= 9)) || ((x == 59) && (y == 5)) || ((x == 60) && (y >= 5 && y <= 9)) ||
              ((x >= 62 && x <= 63) && (y >= 5 && y <= 9)) || ((x == 64) && (y == 5)) || ((x == 64) && (y == 9)) || ((x == 65) && (y >= 5 && y <= 9)) ||
                         
              ((x == 68) && (y == 9)) ||
                         
              ((x == 73) && (y == 6)) || ((x >= 74 && x <= 75) && (y >= 5 && y <= 9)) || ((x == 73) && (y == 9)) || ((x == 76) && (y == 9));

    
    // Display Controls
    wire xrange_3tier_ob = x >= 43 && x <= 53;
    wire xrange_3tier_ib = x >= 47 && x <= 49;
    wire xrange_mid_ib_L = x >= 33 && x <= 35;
    wire xrange_mid_ib_R = x >= 61 && x <= 63;
    wire yrange_top_ob = y >= 18 && y <= 26;
    wire yrange_top_ib = y >= 21 && y <= 23;
    wire yrange_mid_ob = y >= 29 && y <= 37;
    wire yrange_mid_ib = y >= 32 && y <= 34; 
    wire yrange_bottom_ob = y >= 40 && y <= 48;
    wire yrange_bottom_ib = y >= 43 && y <= 45;
    
    wire BUTTONS = ((x == 43) && (yrange_top_ob)) || ((x == 53) && (yrange_top_ob)) || ((xrange_3tier_ob) && (y == 18)) || ((xrange_3tier_ob) && (y == 26)) ||
                   ((x == 45) && (y == 20)) || ((x == 45) && (y == 24)) || ((x == 51) && (y == 20)) || ((x == 51) && (y == 24)) ||
                   ((x == 47) && (yrange_top_ib)) || ((x == 49) && (yrange_top_ib)) || ((xrange_3tier_ib) && (y == 21)) || ((xrange_3tier_ib) && (y == 23)) ||
                   ((x == 48) && (y == 22)) ||      
                   
                   ((x == 43) && (yrange_mid_ob)) || ((x == 53) && (yrange_mid_ob)) || ((xrange_3tier_ob) && (y == 29)) || ((xrange_3tier_ob) && (y == 37)) ||     
                   ((x == 45) && (y == 31)) || ((x == 45) && (y == 35)) || ((x == 51) && (y == 31)) || ((x == 51) && (y == 35)) ||
                   ((x == 47) && (yrange_mid_ib)) || ((x == 49) && (yrange_mid_ib)) || ((xrange_3tier_ib) && (y == 32)) || ((xrange_3tier_ib) && (y == 34)) ||
                   ((x == 48) && (y == 33)) ||
                    
                   ((x == 43) && (yrange_bottom_ob)) || ((x == 53) && (yrange_bottom_ob)) || ((xrange_3tier_ob) && (y == 40)) || ((xrange_3tier_ob) && (y == 48)) ||
                   ((x == 45) && (y == 42)) || ((x == 45) && (y == 46)) || ((x == 51) && (y == 42)) || ((x == 51) && (y == 46)) ||
                   ((x == 47) && (yrange_bottom_ib)) || ((x == 49) && (yrange_bottom_ib)) || ((xrange_3tier_ib) && (y == 43)) || ((xrange_3tier_ib) && (y == 45)) ||      
                   ((x == 48) && (y == 44)) ||
    
                   ((x == 29) && (yrange_mid_ob)) || ((x == 39) && (yrange_mid_ob)) || ((x >= 29 && x <= 39) && (y == 29)) || ((x >= 29 && x <= 39) && (y == 37)) ||     
                   ((x == 31) && (y == 31)) || ((x == 31) && (y == 35)) || ((x == 37) && (y == 31)) || ((x == 37) && (y == 35)) ||
                   ((x == 33) && (yrange_mid_ib)) || ((x == 35) && (yrange_mid_ib)) || ((xrange_mid_ib_L) && (y == 32)) || ((xrange_mid_ib_L) && (y == 34)) ||      
                   ((x == 34) && (y == 33)) ||
    
                   ((x == 57) && (yrange_mid_ob)) || ((x == 67) && (yrange_mid_ob)) || ((x >= 57 && x <= 67) && (y == 29)) || ((x >= 57 && x <= 67) && (y == 37)) ||
                   ((x == 59) && (y == 31)) || ((x == 59) && (y == 35)) || ((x == 65) && (y == 31)) || ((x == 65) && (y == 35)) ||
                   ((x == 61) && (yrange_mid_ib)) || ((x == 63) && (yrange_mid_ib)) || ((xrange_mid_ib_R) && (y == 32)) || ((xrange_mid_ib_R) && (y == 34)) ||
                   ((x == 62) && (y == 33));      
    
    //Display functions
    wire ENTER = ((x == 54) && (y == 38)) || ((x == 55) && (y == 39)) || ((x == 56) && (y == 40)) || ((x == 57) && (y == 41)) || ((x == 58) && (y == 44)) || ((x == 58) && (y == 42)) || 
                 ((x == 59) && (y >= 43 && y <= 44)) || ((x == 60) && (y >= 42 && y <= 44)) ||
    
                 ((x == 61) && (y >= 45 && y <= 49)) || ((x >= 61 && x <= 64) && (y == 45)) || ((x >= 61 && x <= 63) && (y == 47)) || ((x >= 61 && x <= 64) && (y == 49)) ||
                 ((x == 66) && (y >= 45 && y <= 49)) || ((x == 67) && (y == 46)) || ((x == 68) && (y == 47)) || ((x == 69) && (y >= 45 && y <= 49)) ||
                 ((x >= 71 && x <= 75) && (y == 45)) || ((x == 73) && (y >= 45 && y <= 49)) ||
                 ((x == 77) && (y >= 45 && y <= 49)) || ((x >= 77 && x <= 80) && (y == 45)) || ((x >= 77 && x <= 79) && (y == 47)) || ((x >= 77 && x <= 80) && (y == 49)) ||
                 ((x == 82) && (y >= 45 && y <= 49)) || ((x >= 82 && x <= 84) && (y == 45)) || ((x == 85) && (y == 46)) || ((x >= 82 && x <= 84) && (y == 47)) || ((x == 84) && (y == 48)) || ((x == 85) && (y == 49));
    
    wire NEXT = ((x == 62) && (y >= 24 && y <= 28)) || ((x >= 62 && x <= 67) && (y == 24)) || ((x == 68) && (y >= 22 && y <= 26)) || ((x == 69) && (y >= 23 && y <= 25)) || ((x == 70) && (y == 24)) ||
    
                ((x == 72) && (y >= 21 && y <= 25)) || ((x == 73) && (y == 22)) || ((x == 74) && (y == 23)) || ((x == 75) && (y >= 21 && y <= 25)) || 
                ((x == 77) && (y >= 21 && y <= 25)) || ((x >= 77 && x <= 80) && (y == 21)) || ((x >= 77 && x <= 79) && (y == 23)) || ((x >= 77 && x <= 80) && (y == 25)) ||
                ((x == 82) && (y >= 21 && y <= 22)) || ((x == 82) && (y >= 24 && y <= 25)) || ((x >= 83 && x <= 84) && (y == 23)) || ((x == 85) && (y >= 21 && y <= 22)) || ((x == 85) && (y >= 24 && y <= 25)) ||
                ((x >= 87 && x <= 91) && (y == 21)) || ((x == 89) && (y >= 21 && y <= 25));
    
    
    wire GRAB_CHAIR = ((x == 34) && (y >= 24 && y <= 29)) || ((x >= 29 && x <= 34) && (y == 24)) || ((x == 28) && (y >= 22 && y <= 26)) || ((x == 27) && (y >= 23 && y <= 25)) || ((x == 26) && (y == 24)) ||
    
                      ((x >= 6 && x <= 7) && (y == 21)) || ((x == 5) && (y >= 22 && y <= 24)) || ((x >= 6 && x <= 7) && (y == 25)) || ((x == 8) && (y >= 23 && y <= 24)) || ((x == 7) && (y == 23)) ||
                      ((x == 10) && (y >= 21 && y <= 25)) || ((x >= 10 && x <= 12) && (y == 21)) || ((x == 13) && (y == 22)) || ((x >= 11 && x <= 12) && (y == 23)) || ((x == 12) && (y == 24)) || ((x == 13) && (y == 25)) ||
                      ((x == 15) && (y >= 22 && y <= 25)) || ((x >= 16 && x <= 17) && (y == 21)) || ((x >= 15 && x <= 18) && (y == 23)) || ((x == 18) && (y >= 22 && y <= 25)) ||
                      ((x == 20) && (y >= 21 && y <= 25)) || ((x >= 20 && x <= 22) && (y == 21)) || ((x == 23) && (y == 22)) || ((x >= 20 && x <= 22) && (y == 23)) || ((x == 23) && (y == 24)) || ((x >= 20 && x <= 22) && (y == 25)) ||  
    
                      ((x == 8) && (y == 28)) || ((x >= 6 && x <= 7) && (y == 27)) || ((x == 5) && (y >= 28 && y <= 30)) || ((x >= 6 && x <= 7) && (y == 31)) || ((x == 8) && (y == 30)) ||
                      ((x == 10) && (y >= 27 && y <= 31)) || ((x >= 10 && x <= 13) && (y == 29)) || ((x == 13) && (y >= 27 && y <= 31)) ||
                      ((x == 15) && (y >= 28 && y <= 31)) || ((x >= 16 && x <= 17) && (y == 27)) || ((x == 18) && (y >= 28 && y <= 31)) || ((x >= 15 && x <= 18) && (y == 29)) ||
                      ((x >= 20 && x <= 22) && (y == 27)) || ((x == 21) && (y >= 27 && y <= 31)) || ((x >= 20 && x <= 22) && (y == 31)) ||
                      ((x == 24) && (y >= 27 && y <= 31)) || ((x >= 24 && x <= 26) && (y == 27)) || ((x == 27) && (y == 28)) || ((x >= 24 && x <= 26) && (y == 29)) || ((x == 26) && (y == 30)) || ((x == 27) && (y == 31));

    //Display >>>
    wire arrow2 = ((x == 86) && (y == 57)) || ((x == 87) && (y == 58)) || ((x == 86) && (y == 59)) ||
                  ((x == 89) && (y == 57)) || ((x == 90) && (y == 58)) || ((x == 89) && (y == 59)) ||
                  ((x == 92) && (y == 57)) || ((x == 93) && (y == 58)) || ((x == 92) && (y == 59));   

    always @ (*) begin
    oled_data = WHITE;
        if (S1 || BUTTONS || ENTER || NEXT || GRAB_CHAIR) begin
            oled_data = BLACK;
        end
        else if (arrow2) begin
            oled_data = RED;
        end
    end 
endmodule 
