module Game_End_1(
  input [6:0] x,
  input [5:0] y,
  input [8:0] score,
  output reg [15:0] oled_data
);

//Define constant as local parameter
//Colour display
localparam GREEN = 16'h07E0;
localparam ORANGE = 16'hFFE0; //Yellow
localparam RED = 16'hF800;
localparam BLACK = 16'h0000;
localparam PURPLE = 16'hF81F;
localparam YELLOW = 16'hFC00;    
localparam BLUE = 16'h001F;
localparam WHITE = 16'hFFFF;
localparam CYAN = 16'hF81F;
localparam MAGENTA = 16'hF81F;
localparam BROWN = 16'h8204;
localparam SKYBLUE = 16'h5FFF;

wire n1;
wire c;
wire n2;
wire n3;

wire [3:0] num1;
wire [3:0] num2;
wire [3:0] num3;

assign num1 = score / 100;
assign num2 = score % 10;
assign num3 = score % 100;

Number #(.X(3), .Y(3)) number1(x, y, num1, n1);
Colon #(.X(12), .Y(3)) colon(x, y, c);
Number #(.X(18), .Y(3)) number2(x, y, num2, n2);
Number #(.X(27), .Y(3)) number3(x, y, num3, n3);

    //Display Time Taken 
    wire TIME_TAKEN = ((x == 9) && (y == 26)) || ((x == 16) && (y == 26)) || ((x == 15) && (y == 27)) || ((x == 10) && (y >= 25 && y <= 27)) || ((x >= 11 && x <= 12) && (y >= 27 && y <= 30)) || ((x == 14) && (y >= 27 && y <= 30)) ||  ((x >= 10 && x <= 15) && (y == 25)) || ((x == 13) && (y == 31)) ||
                      ((x == 18) && (y == 26)) || ((x == 18) && (y == 30)) || ((x == 23) && (y == 26)) || ((x == 23) && (y == 30)) || ((x == 19) && (y >= 25 && y <= 31)) || ((x == 20) && (y >= 27 && y <= 29)) ||  ((x == 22) && (y >= 27 && y <= 29)) || ((x >= 19 && x <= 22) && (y == 25)) || ((x >= 19 && x <= 22) && (y == 31)) ||
                      ((x == 25) && (y >= 26 && y <= 30)) || ((x == 26) && (y >= 25 && y <= 31)) || ((x == 32) && (y >= 26 && y <= 30)) || ((x == 28) && (y >= 28 && y <= 30)) || ((x == 29) && (y >= 29 && y <= 30)) || ((x == 30) && (y >= 28 && y <= 30)) || ((x == 27) && (y == 25)) || ((x == 27) && (y == 31)) || ((x == 29) && (y == 27)) || ((x == 31) && (y == 31)) ||  ((x >= 28 && x <= 30) && (y == 26)) ||  ((x >= 30 && x <= 31) && (y == 25)) ||
                      ((x == 34) && (y >= 26 && y <= 30)) || ((x == 35) && (y >= 25 && y <= 31)) || ((x >= 35 && x <= 39) && (y == 31)) || ((x >= 35 && x <= 39) && (y == 25)) || ((x >= 37 && x <= 39) && (y == 27)) || ((x >= 37 && x <= 39) && (y == 29)) || ((x == 39) && (y >= 27 && y <= 29)) || ((x == 40) && (y == 26)) || ((x == 40) && (y == 30)) || 
    
                      ((x == 44) && (y == 26)) || ((x == 51) && (y == 26)) || ((x == 45) && (y >= 25 && y <= 27)) || ((x >= 46 && x <= 47) && (y >= 27 && y <= 30)) || ((x == 49) && (y >= 27 && y <= 30)) ||  ((x >= 45 && x <= 50) && (y == 25)) || ((x == 50) && (y == 27)) || ((x == 48) && (y == 31)) ||                  
                      ((x == 53) && (y >= 27 && y <=30)) || ((x == 54) && (y >= 26 && y <= 31)) || ((x == 55) && (y >= 25 && y <= 26)) || ((x == 55) && (y == 31)) || ((x >= 55 && x <= 57) && (y == 25)) || ((x >= 56 && x <= 57) && (y == 27)) || ((x >= 56 && x <= 57) && (y >= 29 && y <= 30)) || ((x == 58) && (y == 26)) || ((x >= 57 && x <= 58) && (y == 31)) || ((x == 59) && (y >= 27 && y <= 30)) || 
                      ((x == 61) && (y >= 26 && y <=30)) || ((x == 62) && (y >= 25 && y <=31)) || ((x == 63) && (y == 25)) || ((x == 63) && (y == 31)) || ((x == 64) && (y >= 26 && y <= 27)) || ((x == 64) && (y >= 29 && y <= 30)) || ((x == 65) && (y >= 25 && y <= 26)) ||  ((x == 65) && (y >= 30 && y <= 31)) || ((x == 66) && (y == 25)) || ((x == 67) && (y == 26)) || ((x == 66) && (y == 27)) || ((x == 65) && (y == 28)) || ((x == 66) && (y == 29)) || ((x == 67) && (y == 30)) || ((x == 66) && (y == 31)) ||
                      ((x == 69) && (y >= 26 && y <= 30)) || ((x == 70) && (y >= 25 && y <= 31)) || ((x >= 70 && x <= 74) && (y == 31)) || ((x >= 70 && x <= 74) && (y == 25)) || ((x >= 72 && x <= 74) && (y == 27)) || ((x >= 72 && x <= 74) && (y == 29)) || ((x == 74) && (y >= 27 && y <= 29)) || ((x == 75) && (y == 26)) || ((x == 75) && (y == 30)) ||                       
                      ((x == 77) && (y >= 26 && y <= 30)) || ((x == 78) && (y >= 25 && y <= 31)) || ((x == 79) && (y == 25)) || ((x == 79) && (y == 31)) || ((x == 80) && (y == 26)) || ((x == 80) && (y >= 28 && y <= 30)) || ((x == 81) && (y >= 25 && y <= 27)) || ((x == 82) && (y == 25)) || ((x == 82) && (y == 31)) || ((x == 81) && (y >= 29 && y <= 30)) || ((x == 83) && (y >= 26 && y <= 30));

    always @ (*) begin
    oled_data = WHITE;
        if (TIME_TAKEN || n1 || c || n2 || n3) begin
            oled_data = BLACK;
        end
    end 

endmodule
