module Game_Screen_1(
  input [6:0] x,
  input [5:0] y,
  output reg [15:0] oled_data
);

//Define constant as local parameter
//Colour display
localparam GREEN = 16'h07E0;
localparam ORANGE = 16'hFFE0; //Yellow
localparam RED = 16'hF800;
localparam BLACK = 16'h0000;
localparam PURPLE = 16'hF81F;
localparam YELLOW = 16'hFC00;    
localparam BLUE = 16'h001F;
localparam WHITE = 16'hFFFF;
localparam CYAN = 16'hF81F;
localparam MAGENTA = 16'hF81F;
localparam BROWN = 16'h8204;
localparam SKYBLUE = 16'h5FFF;

    //Display Wordings on Game Home screen  
    wire FLASHING_CHAIR =((x == 20) && (y >= 28 && y <= 32)) || ((x >= 21 && x <= 23) && (y == 28)) || ((x >= 21 && x <= 22) && (y == 30)) ||
                         ((x == 25) && (y >= 28 && y <= 32)) || ((x >=26 && x <= 28) && (y == 32)) || 
                         ((x == 30) && (y >= 29 && y <= 32)) || ((x >= 31 && x <= 32) && (y == 28)) || ((x >= 31 && x <= 32) && (y == 30)) || ((x == 33) && (y >= 29 && y <= 32)) ||
                         ((x >= 36 && x <= 38) && (y == 28)) || ((x == 35) && (y == 29)) || ((x >= 36 && x <= 37) && (y == 30))  || ((x == 38) && (y == 31)) || ((x >= 35 && x <= 37) && (y == 32)) ||
                         ((x == 40) && (y >= 28 && y <= 32)) || ((x >= 41 && x <= 42) && (y == 30)) || ((x == 43) && (y >= 28 && y <= 32)) ||
                         ((x >= 45 && x <= 47) && (y == 28)) || ((x == 46) && (y >= 28 && y <= 32)) ||
                         ((x == 49) && (y >= 28 && y <= 32)) || ((x == 50) && (y == 29)) || ((x == 51) && (y == 30)) || ((x == 52) && (y >= 28 && y <= 32)) ||
                         ((x == 54) && (y >= 29 && y <= 31)) || ((x >= 55 && x <= 56) && (y == 28)) || ((x >= 55 && x <= 56) && (y == 32)) || ((x == 57) && (y >= 30 && y <= 31)) || ((x == 56) && (y == 30)) ||
                         
                         ((x == 64) && (y == 29)) || ((x >= 62 && x <= 63) && (y == 28)) || ((x == 61) && (y >= 29 && y <= 31)) || ((x >= 62 && x <= 63) && (y == 32)) || ((x == 64) && (y == 31)) ||
                         ((x == 66) && (y >= 28 && y <= 32)) || ((x >= 67 && x <= 68) && (y == 30)) || ((x == 69) && (y >= 28 && y <= 32)) ||
                         ((x == 71) && (y >= 29 && y <= 32)) || ((x >= 72 && x <= 73) && (y == 28)) || ((x == 74) && (y >= 29 && y <= 32)) || ((x >= 72 && x <= 73) && (y == 30)) ||
                         ((x >= 76 && x <= 78) && (y == 28)) || ((x == 77) && (y >= 28 && y <= 32)) || ((x >= 76 && x <= 78) && (y == 32)) ||
                         ((x == 80) && (y >= 28 && y <= 32)) || ((x >= 81 && x <= 82) && (y == 28)) || ((x == 83) && (y == 29)) || ((x >= 81 && x <= 82) && (y == 30)) || ((x == 82) && (y == 31)) || ((x == 83) && (y == 32));
                        
    //Display > Game Control <
    wire GAME_CONTROL = ((x == 18) && (y == 42)) || ((x == 19) && (y == 43)) || ((x == 18) && (y == 44)) ||
                        
                        ((x >= 22 && x <= 23) && (y == 41)) || ((x == 21) && (y >= 42 && y <= 44)) || ((x >= 22 && x <= 23) && (y == 45)) || ((x == 24) && (y >= 43 && y <= 44)) || ((x >= 23 && x <= 24) && (y == 43)) ||
                        ((x >= 27 && x <= 28) && (y == 41)) || ((x == 26) && (y >= 42 && y <= 45)) || ((x >= 26 && x <= 29) && (y == 43)) || ((x == 29) && (y >= 42 && y <= 45)) ||
                        ((x == 31) && (y >= 41 && y <= 45)) || ((x == 32) && (y == 42)) || ((x == 33) && (y == 43)) || ((x == 34) && (y == 42)) || ((x == 35) && (y >= 41 && y <= 45)) ||
                        ((x == 37) && (y >= 41 && y <= 45)) || ((x >= 37 && x <= 40) && (y == 41)) || ((x >= 37 && x <= 39) && (y == 43)) || ((x >= 37 && x <= 40) && (y == 45)) ||
                        
                        ((x == 44) && (y >= 42 && y <= 44)) || ((x >=45 && x <= 46) && (y == 41)) || ((x >= 45 && x <= 46) && (y == 45)) || ((x == 47) && (y == 44)) || ((x == 47) && (y == 42)) ||
                        ((x == 49) && (y >= 42 && y <= 44)) || ((x >= 50 && x <= 51) && (y == 41)) || ((x == 52) && (y >= 42 && y <= 44)) || ((x >= 50 && x <= 51) && (y == 45)) ||
                        ((x == 54) && (y >= 41 && y <= 45)) || ((x == 55) && (y == 42)) || ((x == 56) && (y == 43)) || ((x == 57) && (y >= 41 && y <= 45)) ||
                        ((x >= 59 && x <= 63) && (y == 41)) || ((x == 61) && (y >= 41 && y <= 45)) ||
                        ((x == 65) && (y >= 41 && y <= 45)) || ((x >= 65 && x <= 67) && (y == 41)) || ((x == 68) && (y ==42)) || ((x == 67) && (y == 44)) || ((x >= 65 && x <= 67) && (y == 43)) || ((x == 68) && (y == 45)) ||
                        ((x >= 71 && x <= 72) && (y == 41)) || ((x == 70) && (y >= 42 && y <= 44)) || ((x >= 71 && x <= 72) && (y == 45)) || ((x == 73) && (y >= 42 && y <= 44)) ||
                        ((x == 75) && (y >= 41 && y <= 45)) || ((x >= 75 && x <= 78) && (y == 45)) ||
                        ((x == 81) && (y == 42)) || ((x == 80) && (y == 43)) || ((x == 81) && (y == 44));    

    //Blinking Icon
    wire blink = ((x == 12) && (y == 22)) || ((x == 16) && (y == 22)) ||
                 ((x == 12) && (y == 26)) || ((x == 13) && (y >= 25 && y <= 27)) || ((x == 14) && (y >= 24 && y <= 28)) || ((x == 15) && (y >= 25 && y <= 27)) || ((x == 16) && (y == 26)) ||
                 ((x == 12) && (y == 30)) || ((x == 16) && (y == 30)) ||
                 ((x == 12) && (y == 34)) || ((x == 13) && (y >= 33 && y <= 35)) || ((x == 14) && (y >= 32 && y <= 36)) || ((x == 15) && (y >= 33 && y <= 35)) || ((x == 16) && (y == 34)) ||
                 ((x == 12) && (y == 38)) || ((x == 16) && (y == 38)) ||
                 ((x == 20) && (y == 22)) || ((x == 21) && (y >= 21 && y <= 23)) || ((x == 22) && (y >= 20 && y <= 24)) || ((x == 23) && (y >= 21 && y <= 24)) || ((x == 24) && (y == 22)) ||
                 ((x == 26) && (y == 20)) || ((x == 26) && (y == 24)) ||
                 ((x == 28) && (y == 22)) || ((x == 29) && (y >= 21 && y <= 23)) || ((x == 30) && (y >= 20 && y <= 24)) || ((x == 31) && (y >= 21 && y <= 24)) || ((x == 32) && (y == 22)) ||
                 ((x == 34) && (y == 20)) || ((x == 34) && (y == 24));

    
    //Display >>>
    wire arrow1 = ((x == 86) && (y == 57)) || ((x == 87) && (y == 58)) || ((x == 86) && (y == 59)) ||
                  ((x == 89) && (y == 57)) || ((x == 90) && (y == 58)) || ((x == 89) && (y == 59)) ||
                  ((x == 92) && (y == 57)) || ((x == 93) && (y == 58)) || ((x == 92) && (y == 59));    

endmodule