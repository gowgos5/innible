module Settings(
  input [6:0] x,
  input [5:0] y,
  output reg [15:0] oled_data
);

//Define constant as local parameter
//Colour display
localparam GREEN = 16'h07E0;
localparam ORANGE = 16'hFFE0; //Yellow
localparam RED = 16'hF800;
localparam BLACK = 16'h0000;
localparam PURPLE = 16'hF81F;
localparam YELLOW = 16'hFC00;    
localparam BLUE = 16'h001F;
localparam WHITE = 16'hFFFF;
localparam CYAN = 16'hF81F;
localparam MAGENTA = 16'hF81F;
localparam BROWN = 16'h8204;
localparam SKYBLUE = 16'h5FFF;    

    //Choice
    wire ASK = ((x == 25) && (y >= 9 && y <= 11)) || ((x == 26) && (y >= 8 && y <= 12)) || ((x >= 27 && x <= 28) && (y == 8)) || ((x >= 27 && x <= 28) && (y == 12)) ||
               ((x >= 30 && x <= 31) && (y >= 8 && y <= 12)) || ((x == 32) && (y == 10)) || ((x == 33) && (y >= 8 && y <= 12)) ||
               ((x >= 35 && x <= 36) && (y >= 8 && y <= 12)) || ((x == 37) && (y == 8)) || ((x == 37) && (y == 12)) || ((x == 38) && (y >= 8 && y <= 12)) ||
               ((x >= 40 && x <= 41) && (y >= 8 && y <= 12)) || ((x == 42) && (y == 8)) || ((x == 42) && (y == 12)) || ((x == 43) && (y >= 8 && y <= 12)) ||
               ((x >= 45 && x <= 46) && (y >= 8 && y <= 10)) || ((x >= 47 && x <= 48) && (y >= 10 && y <= 12)) || ((x >= 47 && x <= 48) && (y == 8)) || ((x >= 45 && x <= 46) && (y == 12)) ||
               ((x >= 50 && x <= 51) && (y >= 8 && y <= 12)) || ((x >= 52 && x<= 53) && (y == 8)) || ((x >= 52 && x <= 53) && (y == 12)) || ((x == 52) && (y == 10)) ||
               ((x >= 57 && x <= 58) && (y >= 8 && y <= 12)) || ((x == 59) && (y == 8)) || ((x == 59) && (y == 12)) || ((x == 60) && (y >= 8 && y <= 12)) ||
               ((x >= 62 && x <= 63) && (y >= 8 && y <= 12)) || ((x == 64) && (y == 8)) || ((x == 65) && (y >= 8 && y <= 12)) || 
               ((x >= 67 && x <= 68) && (y >= 8 && y <= 12)) || ((x >= 69 && x <= 70) && (y == 8)) || ((x >= 69 && x <= 70) && (y == 12)) || ((x == 69) && (y == 10)) ||
               
               ((x >= 32 && x <= 33) && (y >= 14 && y <= 16)) || ((x >= 34 && x <= 35) && (y >= 16 && y <= 18)) || ((x >= 34 && x <= 35) && (y == 14)) || ((x >= 32 && x <= 33) && (y == 18)) ||
               ((x >= 37 && x <= 38) && (y >= 14 && y <= 18)) || ((x >= 39 && x <= 40) && (y == 14)) || ((x >= 39 && x <= 40) && (y == 18)) || ((x == 39) && (y == 16)) ||
               ((x >= 42 && x <= 45) && (y == 14)) || ((x >= 43 && x <= 44) && (y >= 14 && y <=18)) ||
               ((x >= 47 && x <= 50) && (y == 14)) || ((x >= 48 && x <= 49) && (y >= 14 && y <= 18)) || 
               ((x >= 52 && x <= 55) && (y == 14)) || ((x >= 52 && x <= 55) && (y == 18)) || ((x >= 53 && x <= 54) && (y >= 14 && y <= 18)) ||
               ((x >= 57 && x <= 58) && (y >= 14 && y <= 18)) || ((x == 59 && y == 14)) || ((x == 60) && (y >= 14 && y <= 18)) || 
               ((x >= 62 && x <= 63) && (y >= 14 && y <= 18)) || ((x >= 64 && x <= 65) && (y == 14)) || ((x == 64) && (y == 18)) || ((x == 65) && (y >= 16 && y <= 18)) || 
               
               ((x >= 45 && x <= 48) && (y == 20)) || ((x >= 46 && x <= 47) && (y >= 20 && y <= 24)) ||
               ((x >= 50 && x <= 51) && (y >= 20 && y <= 24)) || ((x == 52) && (y == 20)) || ((x == 52) && (y == 24)) || ((x == 53) && (y >= 20 && y <= 24)) ||
               
               ((x >= 24 && x <= 25) && (y >= 26 && y <= 30)) || ((x >= 26 && x <= 27) && (y == 26)) || ((x == 26) && (y == 30)) || ((x == 27) && (y >= 28 && y <= 30)) ||
               ((x >= 29 && x <= 30) && (y >= 26 && y <= 30)) || ((x == 31) && (y == 26)) || ((x == 31) && (y == 28)) || ((x == 32) && (y >= 26 && y <= 27)) || ((x == 32) && (y >= 29 && y <= 30)) ||
               ((x >= 34 && x <= 35) && (y >= 26 && y <= 30)) || (( x == 36) && (y == 26)) || ((x == 36) && (y == 28)) || ((x == 37) && (y >= 26 && y <= 30)) ||
               ((x >= 39 && x <= 40) && (y >= 26 && y <= 30)) || ((x == 41) && (y == 26)) || ((x == 41) && (y == 28)) || ((x == 41) && (y == 30)) || ((x == 42) && (y == 27)) || ((x == 42) && (y == 29)) ||
                     
               ((x == 46) && (y >= 27 && y <= 29)) || ((x == 47) && (y >= 26 && y <= 30)) || ((x >= 48 && x <= 49) && (y == 26)) || ((x >= 48 && x <= 49) && (y == 30)) ||
               ((x >= 51 && x <= 52) && (y >= 26 && y <= 30)) || ((x == 53) && (y == 28)) || ((x == 54) && (y >= 26 && y <= 30)) ||
               ((x >= 56 && x <= 57) && (y >= 26 && y <= 30)) || ((x == 58) && (y == 27)) || ((x == 58) && (y == 29)) || ((x == 59) && (y >= 26 && y <= 30)) ||
               ((x >= 61 && x <= 64) && (y == 26)) || ((x >= 61 && x <= 64) && (y == 30)) || ((x >= 62 && x <= 63) && (y >= 26 && y <= 30)) ||
               ((x >= 66 && x <= 67) && (y >= 26 && y <= 30)) || ((x == 68) && (y == 26)) || ((x == 68) && (y == 28)) || ((x == 69) && (y >= 26 && y <= 27)) || ((x == 69) && (y >= 29 && y <= 30));
                     
wire one1 = ((x == 22) && (y == 36)) || ((x >= 23 && x <= 24) && (y >= 35 && y <= 38)) || ((x >= 22 && x <= 25) && (y == 39)) || 
            
            ((x == 30) && (y == 35)) || ((x == 30) && (y == 39)) ||
            
            ((x >= 35 && x <= 36) && (y >= 35 && y <= 39)) || ((x == 37) && (y == 35)) || ((x == 37) && (y == 37)) || ((x == 38) && (y >= 35 && y <= 37)) || 
            ((x >= 40 && x <= 41) && (y >= 35 && y <= 39)) || ((x == 42) && (y == 35)) || ((x == 42) && (y == 37)) || ((x == 43) && (y >= 35 && y <= 36)) || ((x == 43) && (y >= 38 && y <= 39)) ||
            ((x >= 45 && x <= 46) && (y >= 35 && y <= 39))|| ((x >= 47 && x <= 48) && (y == 35)) || ((x == 47) && (y == 37)) || ((x >= 47 && x <= 48) && (y == 39)) ||
            ((x >= 50 && x <= 51) && (y >= 35 && y <= 37)) || ((x >= 52 && x <= 53) && (y >= 37 && y <= 39)) || ((x >= 52 && x <= 53) && (y == 35)) || ((x >= 50 && x <= 51) && (y == 39)) ||
            ((x >= 55 && x <= 56) && (y >= 35 && y <= 37)) || ((x >= 57 && x <= 58) && (y >= 37 && y <= 39)) || ((x >= 57 && x <= 58) && (y == 35)) || ((x >= 55 && x <= 56) && (y == 39)) ||
            
            ((x >= 61 && x <= 62) && (y >= 35 && y <= 38)) || ((x >= 61 && x <= 64) && (y == 39)) || 
            ((x >= 66 && x <= 67) && (y >= 35 && y <= 39))|| ((x >= 68 && x <= 69) && (y == 35)) || ((x == 68) && (y == 37)) || ((x >= 68 && x <= 69) && (y == 39)) ||
            ((x >= 71 && x <= 72) && (y >= 35 && y <= 39))|| ((x >= 73 && x <= 74) && (y == 35)) || ((x == 73) && (y == 37)) ||
            ((x >= 76 && x <= 79) && (y == 35)) || ((x >= 77 && x <= 78) && (y >= 35 && y <= 39));  
            
                     
wire two2 = ((x >= 22 && x <= 24) && (y >= 44 && y <= 45)) || ((x >= 24 && x <= 25) && (y >= 45 && y <= 46)) || ((x >= 22 && x <= 24) && (y >= 47 && y <= 48)) || ((x >= 24 && x <= 25) && (y == 48)) ||
            
            ((x == 30) && (y == 44)) || ((x == 30) && (y == 48)) ||
            
            ((x >= 35 && x <= 36) && (y >= 44 && y <= 48)) || ((x == 37) && (y == 44)) || ((x == 37) && (y == 46)) || ((x == 38) && (y >= 44 && y <= 46)) || 
            ((x >= 40 && x <= 41) && (y >= 44 && y <= 48)) || ((x == 42) && (y == 44)) || ((x == 42) && (y == 46)) || ((x == 43) && (y >= 44 && y <= 45)) || ((x == 43) && (y >= 47 && y <= 48)) ||
            ((x >= 45 && x <= 46) && (y >= 44 && y <= 48))|| ((x >= 47 && x <= 48) && (y == 44)) || ((x == 47) && (y == 46)) || ((x >= 47 && x <= 48) && (y == 48)) ||
            ((x >= 50 && x <= 51) && (y >= 44 && y <= 46)) || ((x >= 52 && x <= 53) && (y >= 46 && y <= 48)) || ((x >= 52 && x <= 53) && (y == 44)) || ((x >= 50 && x <= 51) && (y == 48)) ||
            ((x >= 55 && x <= 56) && (y >= 44 && y <= 46)) || ((x >= 57 && x <= 58) && (y >= 46 && y <= 48)) || ((x >= 57 && x <= 58) && (y == 44)) || ((x >= 55 && x <= 56) && (y == 48)) ||
            
            ((x >= 61 && x <= 62) && (y >= 44 && y <= 48)) || ((x == 63) && (y == 44)) || ((x == 63) && (y == 46)) || ((x == 64) && (y >= 44 && y <= 45)) || ((x == 64) && (y >= 47 && y <= 48)) ||
            ((x >= 66 && x <= 69) && (y == 44)) || ((x >= 67 && x <= 68) && (y >= 45 && y <= 47)) || ((x >= 66 && x <= 69) && (y == 48)) ||
            ((x >= 71 && x <= 72) && (y >= 44 && y <= 48)) || ((x >= 73 && x <= 74) && (y == 44)) || ((x == 73) && (y == 48)) || ((x == 74) && (y >= 46 && y <= 48)) ||
            ((x >= 76 && x <= 77) && (y >= 44 && y <= 48)) || ((x == 78) && (y == 46)) || ((x == 79) && (y >= 44 && y <= 48)) || ((x >= 81 && x <= 84) && (y == 44)) || ((x >= 82 && x <= 83) && (y >= 44 && y <= 48));    
                       
    always @ (*) begin
    oled_data = WHITE;
        if (ASK || one1 || two2) begin
            oled_data = BLACK;
        end
    end  
endmodule
