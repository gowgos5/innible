module Game_End_1(
  input [6:0] x,
  input [5:0] y,
  output reg [15:0] oled_data
);

//Define constant as local parameter
//Colour display
localparam GREEN = 16'h07E0;
localparam ORANGE = 16'hFFE0; //Yellow
localparam RED = 16'hF800;
localparam BLACK = 16'h0000;
localparam PURPLE = 16'hF81F;
localparam YELLOW = 16'hFC00;    
localparam BLUE = 16'h001F;
localparam WHITE = 16'hFFFF;
localparam CYAN = 16'hF81F;
localparam MAGENTA = 16'hF81F;
localparam BROWN = 16'h8204;
localparam SKYBLUE = 16'h5FFF;

    //Display Time Taken 
    wire TIME_TAKEN = ((x == 9) && (y == 26)) || ((x == 16) && (y == 26)) || ((x == 15) && (y == 27)) || ((x == 10) && (y >= 25 && y <= 27)) || ((x >= 11 && x <= 12) && (y >= 27 && y <= 30)) || ((x == 14) && (y >= 27 && y <= 30)) ||  ((x >= 10 && x <= 15) && (y == 25)) || ((x == 13) && (y == 31)) ||
                      ((x == 18) && (y == 26)) || ((x == 18) && (y == 30)) || ((x == 23) && (y == 26)) || ((x == 23) && (y == 30)) || ((x == 19) && (y >= 25 && y <= 31)) || ((x == 20) && (y >= 27 && y <= 29)) ||  ((x == 22) && (y >= 27 && y <= 29)) || ((x >= 19 && x <= 22) && (y == 25)) || ((x >= 19 && x <= 22) && (y == 31)) ||
                      ((x == 25) && (y >= 26 && y <= 30)) || ((x == 26) && (y >= 25 && y <= 31)) || ((x == 32) && (y >= 26 && y <= 30)) || ((x == 28) && (y >= 28 && y <= 30)) || ((x == 29) && (y >= 29 && y <= 30)) || ((x == 30) && (y >= 28 && y <= 30)) || ((x == 27) && (y == 25)) || ((x == 27) && (y == 31)) || ((x == 29) && (y == 27)) || ((x == 31) && (y == 31)) ||  ((x >= 28 && x <= 30) && (y == 26)) ||  ((x >= 30 && x <= 31) && (y == 25)) ||
                      ((x == 34) && (y >= 26 && y <= 30)) || ((x == 35) && (y >= 25 && y <= 31)) || ((x >= 35 && x <= 39) && (y == 31)) || ((x >= 35 && x <= 39) && (y == 25)) || ((x >= 37 && x <= 39) && (y == 27)) || ((x >= 37 && x <= 39) && (y == 29)) || ((x == 39) && (y >= 27 && y <= 29)) || ((x == 40) && (y == 26)) || ((x == 40) && (y == 30)) || 
    
                      ((x == 44) && (y == 26)) || ((x == 51) && (y == 26)) || ((x == 45) && (y >= 25 && y <= 27)) || ((x >= 46 && x <= 47) && (y >= 27 && y <= 30)) || ((x == 49) && (y >= 27 && y <= 30)) ||  ((x >= 45 && x <= 50) && (y == 25)) || ((x == 50) && (y == 27)) || ((x == 48) && (y == 31)) ||                  
                      ((x == 53) && (y >= 27 && y <=30)) || ((x == 54) && (y >= 26 && y <= 31)) || ((x == 55) && (y >= 25 && y <= 26)) || ((x == 55) && (y == 31)) || ((x >= 55 && x <= 57) && (y == 25)) || ((x >= 56 && x <= 57) && (y == 27)) || ((x >= 56 && x <= 57) && (y >= 29 && y <= 30)) || ((x == 58) && (y == 26)) || ((x >= 57 && x <= 58) && (y == 31)) || ((x == 59) && (y >= 27 && y <= 30)) || 
                      ((x == 61) && (y >= 26 && y <=30)) || ((x == 62) && (y >= 25 && y <=31)) || ((x == 63) && (y == 25)) || ((x == 63) && (y == 31)) || ((x == 64) && (y >= 26 && y <= 27)) || ((x == 64) && (y >= 29 && y <= 30)) || ((x == 65) && (y >= 25 && y <= 26)) ||  ((x == 65) && (y >= 30 && y <= 31)) || ((x == 66) && (y == 25)) || ((x == 67) && (y == 26)) || ((x == 66) && (y == 27)) || ((x == 65) && (y == 28)) || ((x == 66) && (y == 29)) || ((x == 67) && (y == 30)) || ((x == 66) && (y == 31)) ||
                      ((x == 69) && (y >= 26 && y <= 30)) || ((x == 70) && (y >= 25 && y <= 31)) || ((x >= 70 && x <= 74) && (y == 31)) || ((x >= 70 && x <= 74) && (y == 25)) || ((x >= 72 && x <= 74) && (y == 27)) || ((x >= 72 && x <= 74) && (y == 29)) || ((x == 74) && (y >= 27 && y <= 29)) || ((x == 75) && (y == 26)) || ((x == 75) && (y == 30)) ||                       
                      ((x == 77) && (y >= 26 && y <= 30)) || ((x == 78) && (y >= 25 && y <= 31)) || ((x == 79) && (y == 25)) || ((x == 79) && (y == 31)) || ((x == 80) && (y == 26)) || ((x == 80) && (y >= 28 && y <= 30)) || ((x == 81) && (y >= 25 && y <= 27)) || ((x == 82) && (y == 25)) || ((x == 82) && (y == 31)) || ((x == 81) && (y >= 29 && y <= 30)) || ((x == 83) && (y >= 26 && y <= 30));

    //Display Best Time
    wire BEST_TIME = ((x == 14) && (y >= 48 && y <= 52)) || ((x == 15) && (y >= 47 && y <= 53)) || ((x >= 15 && x <= 18) && (y == 47)) || ((x == 19) && (y == 48)) || ((x == 20) && (y == 49)) || ((x == 19) && (y == 50)) || ((x == 20) && (y == 51)) || ((x == 19) && (y == 52)) || ((x >= 15 && x <= 18) && (y == 53)) || ((x >= 17 && x <= 18) && (y == 49)) || ((x >= 17 && x <= 18) && (y == 51)) ||
                     ((x == 22) && (y >= 48 && y <= 52)) || ((x == 23) && (y >= 47 && y <= 53)) || ((x >= 23 && x <= 27) && (y == 47)) || ((x >= 23 && x <= 27) && (y == 53)) || ((x >= 25 && x <= 27) && (y == 49)) || ((x >= 25 && x <= 27) && (y == 51)) || ((x == 27) && (y >= 49 && y <= 51)) || ((x == 28) && (y == 48)) || ((x == 28) && (y == 52)) || 
                     ((x >= 32 && x <= 35) && (y == 47)) || ((x == 36) && (y == 48)) || ((x >= 33 && x <= 35) && (y == 49)) || ((x == 35) && (y == 50)) || ((x == 36) && (y == 51)) || ((x == 35) && (y == 52)) || ((x >= 31 && x <= 34) && (y == 53)) || ((x >= 30 && x <= 31) && (y == 52)) || ((x == 31) && (y >= 48 && y <= 53)) || ((x >= 31 && x <= 34) && (y == 51)) || ((x == 32) && (y == 50)) || ((x == 32) && (y >= 47 && y <= 48)) ||                      
                     ((x == 38) && (y == 48)) || ((x == 45) && (y == 48)) || ((x == 39) && (y >= 47 && y <= 49)) || ((x >= 40 && x <= 41) && (y >= 49 && y <= 52)) || ((x == 43) && (y >= 49 && y <= 52)) ||  ((x >= 41 && x <= 42) && (y == 53)) || ((x == 44) && (y == 49)) || ((x >= 39 && x <= 44) && (y == 47)) ||                   

                     ((x == 49) && (y == 48)) || ((x == 56) && (y == 48)) || ((x == 50) && (y >= 47 && y <= 49)) || ((x >= 51 && x <= 52) && (y >= 49 && y <= 52)) || ((x == 54) && (y >= 49 && y <= 52)) ||  ((x >= 52 && x <= 53) && (y == 53)) || ((x == 55) && (y == 49)) || ((x >= 50 && x <= 55) && (y == 47)) ||
                     ((x == 58) && (y == 48)) || ((x == 58) && (y == 52)) || ((x == 63) && (y == 48)) || ((x == 63) && (y == 52)) || ((x == 59) && (y >= 47 && y <= 53)) || ((x == 60) && (y >= 49 && y <= 51)) ||  ((x == 62) && (y >= 49 && y <= 51)) || ((x >= 59 && x <= 62) && (y == 47)) || ((x >= 59 && x <= 62) && (y == 53)) ||
                     ((x == 65) && (y >= 48 && y <= 52)) || ((x == 66) && (y >= 47 && y <= 53)) || ((x == 72) && (y >= 48 && y <= 52)) || ((x == 68) && (y >= 50 && y <= 52)) || ((x == 69) && (y >= 51 && y <= 52)) || ((x == 70) && (y >= 50 && y <= 53)) || ((x == 67) && (y == 47)) || ((x == 67) && (y == 53)) || ((x == 69) && (y == 49)) || ((x == 71) && (y == 53)) ||  ((x >= 68 && x <= 70) && (y == 48)) ||  ((x >= 70 && x <= 71) && (y == 47)) ||
                     ((x == 74) && (y >= 48 && y <= 52)) || ((x == 75) && (y >= 47 && y <= 53)) || ((x >= 75 && x <= 79) && (y == 47)) || ((x >= 75 && x <= 79) && (y == 53)) || ((x >= 77 && x <= 79) && (y == 49)) || ((x >= 77 && x <= 79) && (y == 51)) || ((x == 79) && (y >= 49 && y <= 51)) || ((x == 80) && (y == 48)) || ((x == 80) && (y == 52)); 

    always @ (*) begin
    oled_data = WHITE;
        if (TIME_TAKEN || BEST_TIME) begin
            oled_data = BLACK;
        end
    end 

endmodule
