module Mic_Start(
  input [6:0] x,
  input [5:0] y,
  output reg [15:0] oled_data
);

//Define constant as local parameter
//Colour display
localparam GREEN = 16'h07E0;
localparam ORANGE = 16'hFFE0; //Yellow
localparam RED = 16'hF800;
localparam BLACK = 16'h0000;
localparam PURPLE = 16'hF81F;
localparam YELLOW = 16'hFC00;    
localparam BLUE = 16'h001F;
localparam WHITE = 16'hFFFF;
localparam CYAN = 16'hF81F;
localparam MAGENTA = 16'hF81F;
localparam BROWN = 16'h8204;
localparam SKYBLUE = 16'h5FFF;    
localparam LIGHTGREEN = 16'hAFE5;
localparam DARKGREEN = 16'h632C;
    //Mic Test
    wire MIC_vLine = ((x == 27) && (y >= 34 && y <= 43)) || 
                     ((x == 28) && (y >= 32 && y <= 33)) ||
                     ((x == 29) && (y >= 30 && y <= 31)) || 
                     ((x == 34) && (y >= 26 && y <= 28)) ||
                     ((x >= 36 && x <= 37) && (y >= 30 && y <= 33)) || 
                     ((x == 36) && (y >= 33 && y <= 36)) ||
                     ((x == 35) && (y >= 37 && y <= 43)) ||
                     ((x == 38) && (y >= 26 && y <= 29)) ||
                     ((x == 46) && (y >= 22 && y <= 25));
    
    wire MIC_Body = 
                        ((x >= 30 && x <= 31) && (y == 29)) ||
                        ((x >= 30 && x <= 32) && (y == 31)) ||
                        ((x == 32) && (y == 28)) ||
                        ((x == 33) && (y == 27)) ||
                        ((x >= 33 && x <= 34) && (y == 30)) ||
                        ((x == 35) && (y == 26)) ||
                        ((x >= 35 && x <= 38) && (y == 29)) ||
                        ((x >= 36 && x <= 37) && (y == 25)) ||
                        ((x == 38) && (y == 24)) ||
                        ((x == 39) && (y == 23)) ||
                        ((x >= 39 && x <= 40) && (y == 28)) ||
                        ((x == 40) && (y == 22)) ||
                        ((x == 40) && (y == 24)) ||
                        ((x >= 41 && x <= 45) && (y == 21)) ||
                        ((x == 41) && (y == 25)) ||
                        ((x == 41 && x <= 43) && (y == 27)) ||
                        ((x == 42) && (y == 26)) ||
                        ((x >= 44 && x <= 45) && (y == 26));
        
    //Light Grey
    wire color_Mic_LG = ((x == 30) && (y == 30)) ||
                     ((x == 32) && (y == 29)) ||
                     ((x == 33) && (y == 28)) ||
                     ((x == 38) && (y == 25)) ||
                     ((x == 39) && (y == 24)) ||
                     ((x == 39) && (y == 27)) ||
                     ((x == 40) && (y == 26)) ||
                     ((x == 41) && (y == 23)) ||
                     ((x == 42) && (y == 22)) ||
                     ((x == 43) && (y == 26)) ||
                     ((x == 44) && (y == 25)) ||
                     ((x == 44) && (y == 22)) ||
                     ((x == 45) && (y == 22)) ||              
                     ((x == 45) && (y == 23));
    
    //Dark Grey
    wire color_Mic_DG = ((x >= 31 && x <= 32) && (y == 30)) ||
                        ((x >= 33 && x <= 34) && (y == 29)) ||
                        ((x == 35) && (y >= 27 && y <= 28)) ||
                        ((x >= 36 && x <= 37) && (y >= 26 && y <= 28)) ||
                        ((x == 39) && (y >= 25 && y <= 26)) ||
                        ((x == 40) && (y == 25)) ||
                        ((x == 40) && (y == 27)) ||
                        ((x == 41) && (y == 26)) ||
                        ((x == 40) && (y == 23)) || 
                        ((x == 41) && (y == 22)) ||
                        ((x == 43) && (y == 22)) ||
                        ((x == 44) && (y >= 23 && y <= 24)) ||
                        ((x == 45) && (y >= 24 && y <= 25)) ||              
                        ((x >= 42 && x <= 43) && (y >= 23 && y <= 25)) ||                 
                        ((x == 41) && (y == 24));
      
    wire MIC_TEST = ((x == 47) && (y >= 30 && y <= 34)) || ((x == 48) && (y >= 29 && y <= 35)) || ((x == 49) && (y == 29)) || ((x == 49) && (y == 35)) || ((x == 51) && (y == 31)) || ((x == 50) && (y == 32)) || ((x == 52) && (y == 32)) || ((x >= 50 && x <= 52) && (y == 30)) || ((x >= 50 && x <= 52) && (y >= 33 && y <= 34)) || ((x == 53) && (y == 35)) || ((x >= 52 && x <= 53) && (y == 29)) || ((x == 54) && (y >= 30 && y <= 34)) ||
                    ((x == 56) && (y == 56)) || ((x == 56) && (y == 34)) || ((x == 57) && (y >= 29 && y <= 35)) || ((x == 58) && (y >= 31 && y <= 33)) || ((x == 60) && (y >= 31 && y <= 33)) || ((x >= 58 && x <= 60) && (y == 29)) || ((x >= 58 && x <= 60) && (y == 35)) || ((x == 61) && (y == 30)) || ((x == 61) && (y == 34)) ||
                    ((x == 63) && (y >= 31 && y <= 33))  || ((x == 64) && (y >= 30 && y <= 34)) || ((x == 65) && (y >= 29 && y <= 30)) || ((x == 65) && (y >= 34 && y <= 35)) || ((x >= 66 && x <= 67) && (y == 29)) || ((x >= 66 && x <= 67) && (y ==35)) || ((x == 68) && (y == 30)) || ((x == 68) && (y == 34)) || ((x == 66) && (y >= 31 && y <= 33)) || ((x == 67) && (y == 31)) || ((x == 67) && (y == 33)) ||
                    
                    ((x == 47) && (y == 38)) || ((x == 48) && (y >= 37 && y <= 39)) || ((x >= 49 && x <= 53) && (y == 37)) || ((x == 54) && (y == 38)) || ((x == 53) && (y == 39)) || ((x == 52) && (y >= 39 && y <= 42)) || ((x == 51) && (y == 43)) || ((x >= 49 && x <= 50) && (y >= 39 && y <= 42)) ||
                    ((x == 56) && (y >= 38 && y <= 42)) || ((x == 57) && (y >= 37 && y <= 43)) || ((x >= 58 && x <= 61) && (y == 37)) || ((x >= 58 && x <= 61) && (y == 43)) || ((x == 62) && (y == 38)) || ((x == 62) && (y == 42)) || ((x == 61) && (y >= 39 && y <= 41)) || ((x >= 59 && x <= 60) && (y == 39)) || ((x >= 59 && x <= 60) && (y == 41)) ||
                    ((x == 64) && (y == 39)) || ((x == 64) && (y == 42)) || ((x == 65) && (y >= 38 && y <= 43)) || ((x == 66) && (y == 38)) || ((x >= 66 && x <= 69) && (y == 37)) || ((x == 70) && (y == 38)) || ((x >=67 && x <= 69) && (y == 39)) || ((x == 69) && (y == 40)) || ((x == 70) && (y == 41)) || ((x == 69) && (y == 42)) || ((x >= 66 && x <= 68) && (y == 43)) || ((x >= 66 && x <= 68) && (y == 41)) || ((x == 66) && (y == 40)) ||
                    ((x == 72) && (y == 38)) || ((x == 73) && (y >= 37 && y <= 39)) || ((x >= 74 && x <= 78) && (y == 37)) || ((x == 79) && (y == 38)) || ((x == 78) && (y == 39)) || ((x == 77) && (y >= 39 && y <= 42)) || ((x == 76) && (y == 43)) || ((x >= 74 && x <= 75) && (y >= 40 && y <= 42));   
    
    always @ (*) begin
    oled_data = WHITE;
        if (MIC_vLine || MIC_TEST || MIC_Body) begin
            oled_data = BLACK;
        end
        else if (color_Mic_LG) begin
            oled_data = LIGHTGREEN;
        end
        else if (color_Mic_DG) begin
            oled_data = DARKGREEN;
        end
    end  


endmodule

