module Game_Screen_8(
  input [6:0] x,
  input [5:0] y,
  output reg [15:0] oled_data
);

//Define constant as local parameter
//Colour display
localparam GREEN = 16'h07E0;
localparam ORANGE = 16'hFFE0; //Yellow
localparam RED = 16'hF800;
localparam BLACK = 16'h0000;
localparam PURPLE = 16'hF81F;
localparam YELLOW = 16'hFC00;    
localparam BLUE = 16'h001F;
localparam WHITE = 16'hFFFF;
localparam CYAN = 16'hF81F;
localparam MAGENTA = 16'hF81F;
localparam BROWN = 16'h8204;
localparam SKYBLUE = 16'h5FFF;
localparam LIGHTGREEN = 16'hAFE5;

    //Display Loading Game
    wire LOADING_GAME = ((x == 10) && (y >= 17 && y <= 21)) || ((x >= 10 && x <= 13) && (y == 21)) ||
                        ((x == 15) && (y >= 18 && y <= 20)) || ((x >= 16 && x <= 17) && (y == 17)) || ((x == 18) && (y >= 18 && y <= 20)) || ((x >= 16 && x <= 17) && (y == 21)) ||
                        ((x == 20) && (y >= 18 && y <= 21)) || ((x >= 21 && x <= 22) && (y == 17)) || ((x >= 20 && x <= 23) && (y == 19)) || ((x == 23) && (y >= 18 && y <= 21)) ||
                        ((x == 25) && (y >= 17 && y <= 21)) || ((x >= 25 && x <= 27) && (y == 17)) ||  ((x >= 25 && x <= 27) && (y == 21)) || ((x == 28) && (y >= 18 && y <= 20)) ||
                        ((x >= 30 && x <= 32) && (y == 17)) || ((x == 31) && (y >= 17 && y <= 21)) || ((x >= 30 && x <= 32) && (y == 21)) ||
                        ((x == 34) && (y >= 17 && y <= 21)) || ((x == 35) && (y == 18)) || ((x == 36) && (y == 19)) || ((x == 37) && (y >= 17 && y <= 21)) ||
                        ((x == 39) && (y >= 18 && y <= 20)) || ((x >= 40 && x <= 41) && (y == 17)) || ((x >= 40 && x <= 41) && (y == 21)) || ((x == 42) && (y >= 19 && y <= 20)) || ((x >= 41 && x <= 42) && (y == 19)) ||  
    
                        ((x == 46) && (y >= 18 && y <= 20)) || ((x >= 47 && x <= 48) && (y == 17)) || ((x >= 47 && x <= 48) && (y == 21)) || ((x == 49) && (y >= 19 && y <= 20)) || ((x >= 48 && x <= 49) && (y == 19)) ||  
                        ((x == 51) && (y >= 18 && y <= 21)) || ((x >= 52 && x <= 53) && (y == 17)) || ((x >= 51 && x <= 54) && (y == 19)) || ((x == 54) && (y >= 18 && y <= 21)) ||
                        ((x == 56) && (y >= 17 && y <= 21)) || ((x == 57) && (y == 18)) || ((x == 58) && (y == 19)) || ((x == 59) && (y == 18)) || ((x == 60) && (y >= 17 && y <= 21)) ||
                        ((x == 62) && (y >= 17 && y <= 21)) || ((x >= 62 && x <= 65) && (y == 17)) || ((x >= 62 && x <= 64) && (y == 19)) || ((x >= 62 && x <= 65) && (y == 21));
    
    wire LOADING_BAR_OB = ((x >= 10 && x <= 12) && (y >= 29 && y <= 46)) || ((x >= 87 && x <= 89) && (y >= 29 && y <= 46)) ||
                          ((x >= 13 && x <= 86) && (y >= 26 && y <= 28)) || ((x >= 13 && x <= 86) && (y >= 47 && y <= 49));
                          
    wire LOADING_BAR = ((x >= 14 && x <= 30) && (y >= 30 && y <= 45)) ||
                       ((x >= 32 && x <= 49) && (y >= 30 && y <= 45)) ||
                       ((x >= 51 && x <= 67) && (y >= 30 && y <= 45)) ||
                       ((x >= 69 && x <= 85) && (y >= 30 && y <= 45));
    
    wire rule =  ((x >= 12 && x <= 13) && (y == 51)) || ((x >= 10 && x <= 11) && (y >= 51 && y <= 55)) || ((x >= 12 && x <= 13) && (y == 55)) || ((x == 13) && (y >= 53 && y <= 55)) ||
                 ((x >= 15 && x <= 16) && (y >= 51 && y <= 55)) || ((x == 17) && (y == 51)) || ((x == 17 ) && (y == 53)) || ((x == 18) && (y >= 51 && y <= 52)) || ((x == 18) && (y >= 54 && y <= 55)) ||
                 ((x >= 20 && x <= 21) && (y >= 51 && y <= 55)) || ((x == 22) && (y == 51)) || ((x == 22 ) && (y == 53)) || ((x == 23) && (y >= 51 && y <= 55)) ||
                 ((x >= 25 && x <= 26) && (y >= 51 && y <= 55)) || ((x == 27) && (y == 51)) || ((x == 27 ) && (y == 53)) || ((x == 27 ) && (y == 55)) || ((x == 28 ) && (y == 52)) || ((x == 28) && (y == 54)) ||
                     
                 ((x >= 32 && x <= 35) && (y == 51)) || ((x >= 33 && x <= 34) && (y >= 51 && y <= 55)) ||
                 ((x >= 37 && x <= 38) && (y >= 51 && y <= 55)) || ((x == 39) && (y == 53)) || ((x == 40) && (y >= 51 && y <= 55)) || 
                 ((x >= 42 && x <= 43) && (y >= 51 && y <= 55)) || ((x == 44) && (y == 53)) || ((x >= 44 && x <= 45) && (y == 51)) || ((x >= 44 && x <= 45) && (y == 55)) || 
                     
                 ((x == 49) && (y >= 52 && y <= 54)) || ((x == 50) && (y >= 51 && y <= 55)) || ((x >= 51 && x <= 52) && (y == 51)) || ((x >= 51 && x <= 52) && (y == 55)) || 
                 ((x >= 54 && x <= 55) && (y >= 51 && y <= 55)) || ((x == 56) && (y == 53)) || ((x == 57 )&& (y >= 51 && y <= 55)) ||
                 ((x >= 59 && x <= 60) && (y >= 51 && y <= 55)) || ((x == 61) && (y == 51)) || ((x == 61 ) && (y == 53)) || ((x == 62) && (y >= 51 && y <= 55)) ||
                 ((x >= 64 && x <= 67) && (y == 51)) || ((x >= 64 && x <= 67) && (y == 55)) || ((x >= 65 && x <= 66) && (y >= 51 && y < 55)) || 
                 ((x >= 69 && x <= 70) && (y >= 51 && y <= 55)) || ((x == 71 ) && (y == 51)) || ((x == 71 ) && (y == 53)) || ((x == 72) && (y >= 51 && y <= 52)) || ((x == 72) && (y >= 54 && y <= 55)) ||     
                     
                 ((x >= 76 && x <= 77) && (y >= 51 && y <= 55)) || ((x == 78 ) && (y == 51)) || ((x == 78 ) && (y == 53)) || ((x == 78 ) && (y == 55)) || ((x == 79 ) && (y == 52)) || ((x == 79) && (y == 54)) ||
                 ((x == 81) && (y >= 51 && y <= 53)) || ((x == 82) && (y == 53)) || ((x >= 83 && x <= 84) && (y >= 51 && y <= 55)) ||
                 
                 ((x >= 10 && x <= 13) && (y == 57)) || ((x >= 10 && x <= 13) && (y == 61)) || ((x >= 11 && x <= 12) && (y >= 57 && y <= 61)) ||
                 ((x >= 15 && x <= 18) && (y == 57)) || ((x >= 16 && x <= 17) && (y >= 57 && y <= 61)) ||
                 
                 ((x >= 22 && x <= 23) && (y >= 57 && y <= 59)) || ((x >= 24 && x <= 25) && (y == 57)) || ((x >= 24 && x <= 25) && (y >= 59 && y <= 61)) || ((x >= 22 && x <= 23) && (y == 61)) ||
                 ((x >= 27 && x <= 30) && (y == 57)) || ((x >= 28 && x <= 29) && (y >= 57 && y <= 61)) || 
                 ((x >= 32 && x <= 33) && (y >= 57 && y <= 61)) || ((x == 34) && (y == 57)) || ((x == 34) && (y == 61)) || ((x == 35) && (y >= 57 && y <= 61)) || 
                 ((x >= 37 && x <= 38) && (y >= 57 && y <= 61)) || ((x == 39) && (y == 57)) || ((x == 39) && (y == 59)) || ((x == 40) && (y >= 57 && y <= 59)) ||
                 ((x >= 42 && x <= 43) && (y >= 57 && y <= 59)) || ((x >= 44 && x <= 45) && (y == 57)) || ((x >= 44 && x <= 45) && (y >= 59 && y <= 61)) || ((x >= 42 && x <= 43) && (y == 61)) ||

                 ((x >= 49 && x <= 50) && (y >= 57 && y <= 61)) || ((x >= 51 && x <= 52) && (y == 57)) || ((x == 51) && (y == 59)) ||
                 ((x >= 54 && x <= 55) && (y >= 57 && y <= 61)) || ((x >= 56 && x <= 57) && (y == 61)) ||
                 ((x >= 59 && x <= 60) && (y >= 57 && y <= 61)) || ((x == 61) && (y == 57)) || ((x == 61) && (y == 59)) || ((x == 62) && (y >= 57 && y <= 61)) ||
                 ((x >= 64 && x <= 65) && (y >= 57 && y <= 59)) || ((x >= 66 && x <= 67) && (y == 57)) || ((x >= 66 && x <= 67) && (y >= 59 && y <= 61)) || ((x >= 64 && x <= 65) && (y == 61)) ||
                 ((x >= 69 && x <= 70) && (y >= 57 && y <= 61)) || ((x == 71) && (y == 59)) || ((x == 72) && (y >= 57 && y <= 61)) || 
                 ((x >= 74 && x <= 77) && (y == 57)) || ((x >= 74 && x <= 77) && (y == 61)) || ((x >= 75 && x <= 76) && (y >= 57 && y <= 61)) ||
                 ((x >= 79 && x <= 80) && (y >= 57 && y <= 61)) || ((x == 81) && (y == 57)) || ((x == 82) && (y >= 57 && y <= 61)) ||
                 ((x >= 84 && x <= 85) && (y >= 57 && y <= 61)) || ((x == 86) && (y == 57)) || ((x == 86) && (y == 61)) || ((x == 87) && (y == 57)) || ((x == 87) && (y >= 59 && y <= 61));

    always @ (*) begin
    oled_data = WHITE;
        if (LOADING_GAME || LOADING_BAR_OB) begin
            oled_data = BLACK;
        end
        else if (LOADING_BAR) begin
            oled_data = LIGHTGREEN; 
        end
        else if (rule) begin
            oled_data = RED;
        end
    end 

endmodule

